module imem (
	input  [ 5:0] addr,
	output reg [31:0] data
);

	// echo -e {00..63}": data = 32'h00000000;\n"
	// xx : data = {6'dx,5'dx,5'dx,5'dx,5'dx,6'dx};
	always @(addr) begin
		case(addr)
			00 : data = 32'h00001820;
			01 : data = 32'h2001000A;
			02 : data = 32'h00231820;
			03 : data = 32'hAC030001;
			04 : data = 32'h28210001;
			05 : data = 32'h00012029;
			06 : data = 32'h1480fff6;
			07 : data = 32'h8C030001;
			08 : data = 32'h00000000;
			09 : data = 32'h00000000;
			10 : data = 32'h00000000;
			11 : data = 32'h00000000;
			12 : data = 32'h00000000;
			13 : data = 32'h00000000;
			14 : data = 32'h00000000;
			15 : data = 32'h00000000;
			16 : data = 32'h00000000;
			17 : data = 32'h00000000;
			18 : data = 32'h00000000;
			19 : data = 32'h00000000;
			20 : data = 32'h00000000;
			21 : data = 32'h00000000;
			22 : data = 32'h00000000;
			23 : data = 32'h00000000;
			24 : data = 32'h00000000;
			25 : data = 32'h00000000;
			26 : data = 32'h00000000;
			27 : data = 32'h00000000;
			28 : data = 32'h00000000;
			29 : data = 32'h00000000;
			30 : data = 32'h00000000;
			31 : data = 32'h00000000;
			32 : data = 32'h00000000;
			33 : data = 32'h00000000;
			34 : data = 32'h00000000;
			35 : data = 32'h00000000;
			36 : data = 32'h00000000;
			37 : data = 32'h00000000;
			38 : data = 32'h00000000;
			39 : data = 32'h00000000;
			40 : data = 32'h00000000;
			41 : data = 32'h00000000;
			42 : data = 32'h00000000;
			43 : data = 32'h00000000;
			44 : data = 32'h00000000;
			45 : data = 32'h00000000;
			46 : data = 32'h00000000;
			47 : data = 32'h00000000;
			48 : data = 32'h00000000;
			49 : data = 32'h00000000;
			50 : data = 32'h00000000;
			51 : data = 32'h00000000;
			52 : data = 32'h00000000;
			53 : data = 32'h00000000;
			54 : data = 32'h00000000;
			55 : data = 32'h00000000;
			56 : data = 32'h00000000;
			57 : data = 32'h00000000;
			58 : data = 32'h00000000;
			59 : data = 32'h00000000;
			60 : data = 32'h00000000;
			61 : data = 32'h00000000;
			62 : data = 32'h00000000;
			63 : data = 32'h00000000;
		endcase
	end

endmodule
